package const_MEM is

   constant ADDRESS_LENGTH_IN : natural := 32; -- input address length
   constant ADDRESS_LENGTH : natural := 8; -- effective address length to avoid overflow
   constant DATA_LENGTH : natural := 32;

end const_MEM;