package alu_types is
	type TYPE_OP is (ADD, SUB, MULT, BITAND, BITOR, BITXOR, FUNCSLT, FUNCLSL, FUNCLSR, FUNCRL, FUNCRR);
end alu_types;
