library verilog;
use verilog.vl_types.all;
entity tb_iir_LA is
end tb_iir_LA;
