library IEEE;
use IEEE.std_logic_1164.all;

entity Mult_Dadda32 is
	generic( N : natural := 32);
	port( x : in std_logic_vector(N - 1 downto 0);
		y : in std_logic_vector(N - 1 downto 0);
		z : out std_logic_vector(2*N - 1 downto 0));
end entity Mult_Dadda32;

architecture arch of Mult_Dadda32 is
component full_adder is
	port(
		a : in std_logic;
		b : in std_logic;
		cin : in  std_logic;
		s : out std_logic;
		cout : out std_logic);
end component;

component half_adder is
	port(
		a : in std_logic;
		b : in std_logic;
		s : out std_logic;
		cout : out std_logic);
end component;

component mbe_ppst is
	generic(n : natural := 32);
	port(triplet : in std_logic_vector(2 downto 0);--sign bit representation
		Y : in std_logic_vector(N-1 downto 0);
		pp : out std_logic_vector(N downto 0);
		S : out std_logic);
end component;

type P_t is array (N/2 downto 0) of std_logic_vector(N downto 0);
signal P : P_t;
signal Sig, nSig : std_logic_vector(N/2 downto 0);
subtype Sum_t is std_logic_vector(588 downto 0);
signal Sum : Sum_t;
subtype Cout_t is std_logic_vector(588 downto 0);
signal Cout : Cout_t;
signal ppg0_three_digits, ppglast_three_digits : std_logic_vector(2 downto 0);

begin

ppg0_three_digits <= x(1 downto 0)&'0';
ppg0: mbe_ppst generic map(N) port map(ppg0_three_digits, y, P(0), Sig(0));

F0: for i in 1 to n/2-1 generate
	ppgi: mbe_ppst generic map(N) port map(x((2*i + 1) downto (2*i - 1)), y, P(i), Sig(i));
end generate;

ppglast_three_digits(N - 2*(N/2) downto 0) <= x(n - 1 downto 2*(n/2) -1);ppglast_three_digits(2 downto N - 2*(N/2) + 1) <= (others => '0');
ppglast: mbe_ppst generic map(N) port map(ppglast_three_digits, y, P(n/2), Sig(n/2));

HA1 : half_adder port map(Sig(12), P(12)(0), Sum(0), Cout(0));
HA2 : half_adder port map(P(12)(1), P(11)(3), Sum(1), Cout(1));
FA1 : full_adder port map(Sig(13), P(13)(0), P(12)(2), Sum(2), Cout(2));
HA3 : half_adder port map(P(11)(4), P(10)(6), Sum(3), Cout(3));
FA2 : full_adder port map(P(13)(1), P(12)(3), P(11)(5), Sum(4), Cout(4));
HA4 : half_adder port map(P(10)(7), P(9)(9), Sum(5), Cout(5));
FA3 : full_adder port map(Sig(14), P(14)(0), P(13)(2), Sum(6), Cout(6));
FA4 : full_adder port map(P(12)(4), P(11)(6), P(10)(8), Sum(7), Cout(7));
HA5 : half_adder port map(P(9)(10), P(8)(12), Sum(8), Cout(8));
FA5 : full_adder port map(P(14)(1), P(13)(3), P(12)(5), Sum(9), Cout(9));
FA6 : full_adder port map(P(11)(7), P(10)(9), P(9)(11), Sum(10), Cout(10));
HA6 : half_adder port map(P(8)(13), P(7)(15), Sum(11), Cout(11));
FA7 : full_adder port map(Sig(15), P(15)(0), P(14)(2), Sum(12), Cout(12));
FA8 : full_adder port map(P(13)(4), P(12)(6), P(11)(8), Sum(13), Cout(13));
FA9 : full_adder port map(P(10)(10), P(9)(12), P(8)(14), Sum(14), Cout(14));
HA7 : half_adder port map(P(7)(16), P(6)(18), Sum(15), Cout(15));
FA10 : full_adder port map(P(15)(1), P(14)(3), P(13)(5), Sum(16), Cout(16));
FA11 : full_adder port map(P(12)(7), P(11)(9), P(10)(11), Sum(17), Cout(17));
FA12 : full_adder port map(P(9)(13), P(8)(15), P(7)(17), Sum(18), Cout(18));
HA8 : half_adder port map(P(6)(19), P(5)(21), Sum(19), Cout(19));
FA13 : full_adder port map(P(16)(0), P(15)(2), P(14)(4), Sum(20), Cout(20));
FA14 : full_adder port map(P(13)(6), P(12)(8), P(11)(10), Sum(21), Cout(21));
FA15 : full_adder port map(P(10)(12), P(9)(14), P(8)(16), Sum(22), Cout(22));
FA16 : full_adder port map(P(7)(18), P(6)(20), P(5)(22), Sum(23), Cout(23));
FA17 : full_adder port map(Sig(0), P(1)(31), P(2)(29), Sum(24), Cout(24));
FA18 : full_adder port map(P(3)(27), P(4)(25), P(5)(23), Sum(25), Cout(25));
FA19 : full_adder port map(P(6)(21), P(7)(19), P(8)(17), Sum(26), Cout(26));
FA20 : full_adder port map(P(9)(15), P(10)(13), P(11)(11), Sum(27), Cout(27));
FA21 : full_adder port map(Sig(0), P(1)(32), P(2)(30), Sum(28), Cout(28));
FA22 : full_adder port map(P(3)(28), P(4)(26), P(5)(24), Sum(29), Cout(29));
FA23 : full_adder port map(P(6)(22), P(7)(20), P(8)(18), Sum(30), Cout(30));
FA24 : full_adder port map(P(9)(16), P(10)(14), P(11)(12), Sum(31), Cout(31));
FA25 : full_adder port map(nSig(0), nSig(1), P(2)(31), Sum(32), Cout(32));
FA26 : full_adder port map(P(3)(29), P(4)(27), P(5)(25), Sum(33), Cout(33));
FA27 : full_adder port map(P(6)(23), P(7)(21), P(8)(19), Sum(34), Cout(34));
FA28 : full_adder port map(P(9)(17), P(10)(15), P(11)(13), Sum(35), Cout(35));
FA29 : full_adder port map('1', P(2)(32), P(3)(30), Sum(36), Cout(36));
FA30 : full_adder port map(P(4)(28), P(5)(26), P(6)(24), Sum(37), Cout(37));
FA31 : full_adder port map(P(7)(22), P(8)(20), P(9)(18), Sum(38), Cout(38));
HA9 : half_adder port map(P(10)(16), P(11)(14), Sum(39), Cout(39));
FA32 : full_adder port map(nSig(2), P(3)(31), P(4)(29), Sum(40), Cout(40));
FA33 : full_adder port map(P(5)(27), P(6)(25), P(7)(23), Sum(41), Cout(41));
FA34 : full_adder port map(P(8)(21), P(9)(19), P(10)(17), Sum(42), Cout(42));
FA35 : full_adder port map('1', P(3)(32), P(4)(30), Sum(43), Cout(43));
FA36 : full_adder port map(P(5)(28), P(6)(26), P(7)(24), Sum(44), Cout(44));
HA10 : half_adder port map(P(8)(22), P(9)(20), Sum(45), Cout(45));
FA37 : full_adder port map(nSig(3), P(4)(31), P(5)(29), Sum(46), Cout(46));
FA38 : full_adder port map(P(6)(27), P(7)(25), P(8)(23), Sum(47), Cout(47));
FA39 : full_adder port map('1', P(4)(32), P(5)(30), Sum(48), Cout(48));
HA11 : half_adder port map(P(6)(28), P(7)(26), Sum(49), Cout(49));
FA40 : full_adder port map(nSig(4), P(5)(31), P(6)(29), Sum(50), Cout(50));
HA12 : half_adder port map('1', P(5)(32), Sum(51), Cout(51));
HA13 : half_adder port map(Sig(8), P(8)(0), Sum(52), Cout(52));
HA14 : half_adder port map(P(8)(1), P(7)(3), Sum(53), Cout(53));
FA41 : full_adder port map(Sig(9), P(9)(0), P(8)(2), Sum(54), Cout(54));
HA15 : half_adder port map(P(7)(4), P(6)(6), Sum(55), Cout(55));
FA42 : full_adder port map(P(9)(1), P(8)(3), P(7)(5), Sum(56), Cout(56));
HA16 : half_adder port map(P(6)(7), P(5)(9), Sum(57), Cout(57));
FA43 : full_adder port map(Sig(10), P(10)(0), P(9)(2), Sum(58), Cout(58));
FA44 : full_adder port map(P(8)(4), P(7)(6), P(6)(8), Sum(59), Cout(59));
HA17 : half_adder port map(P(5)(10), P(4)(12), Sum(60), Cout(60));
FA45 : full_adder port map(P(10)(1), P(9)(3), P(8)(5), Sum(61), Cout(61));
FA46 : full_adder port map(P(7)(7), P(6)(9), P(5)(11), Sum(62), Cout(62));
HA18 : half_adder port map(P(4)(13), P(3)(15), Sum(63), Cout(63));
FA47 : full_adder port map(Sig(11), P(11)(0), P(10)(2), Sum(64), Cout(64));
FA48 : full_adder port map(P(9)(4), P(8)(6), P(7)(8), Sum(65), Cout(65));
FA49 : full_adder port map(P(6)(10), P(5)(12), P(4)(14), Sum(66), Cout(66));
HA19 : half_adder port map(P(3)(16), P(2)(18), Sum(67), Cout(67));
FA50 : full_adder port map(P(11)(1), P(10)(3), P(9)(5), Sum(68), Cout(68));
FA51 : full_adder port map(P(8)(7), P(7)(9), P(6)(11), Sum(69), Cout(69));
FA52 : full_adder port map(P(5)(13), P(4)(15), P(3)(17), Sum(70), Cout(70));
HA20 : half_adder port map(P(2)(19), P(1)(21), Sum(71), Cout(71));
FA53 : full_adder port map(P(11)(2), P(10)(4), P(9)(6), Sum(72), Cout(72));
FA54 : full_adder port map(P(8)(8), P(7)(10), P(6)(12), Sum(73), Cout(73));
FA55 : full_adder port map(P(5)(14), P(4)(16), P(3)(18), Sum(74), Cout(74));
FA56 : full_adder port map(P(2)(20), P(1)(22), P(0)(24), Sum(75), Cout(75));
FA57 : full_adder port map(P(10)(5), P(9)(7), P(8)(9), Sum(76), Cout(76));
FA58 : full_adder port map(P(7)(11), P(6)(13), P(5)(15), Sum(77), Cout(77));
FA59 : full_adder port map(P(4)(17), P(3)(19), P(2)(21), Sum(78), Cout(78));
FA60 : full_adder port map(P(1)(23), P(0)(25), Cout(0), Sum(79), Cout(79));
FA61 : full_adder port map(P(9)(8), P(8)(10), P(7)(12), Sum(80), Cout(80));
FA62 : full_adder port map(P(6)(14), P(5)(16), P(4)(18), Sum(81), Cout(81));
FA63 : full_adder port map(P(3)(20), P(2)(22), P(1)(24), Sum(82), Cout(82));
FA64 : full_adder port map(P(0)(26), Cout(1), Sum(2), Sum(83), Cout(83));
FA65 : full_adder port map(P(8)(11), P(7)(13), P(6)(15), Sum(84), Cout(84));
FA66 : full_adder port map(P(5)(17), P(4)(19), P(3)(21), Sum(85), Cout(85));
FA67 : full_adder port map(P(2)(23), P(1)(25), P(0)(27), Sum(86), Cout(86));
FA68 : full_adder port map(Cout(2), Cout(3), Sum(4), Sum(87), Cout(87));
FA69 : full_adder port map(P(7)(14), P(6)(16), P(5)(18), Sum(88), Cout(88));
FA70 : full_adder port map(P(4)(20), P(3)(22), P(2)(24), Sum(89), Cout(89));
FA71 : full_adder port map(P(1)(26), P(0)(28), Cout(4), Sum(90), Cout(90));
FA72 : full_adder port map(Cout(5), Sum(6), Sum(7), Sum(91), Cout(91));
FA73 : full_adder port map(P(6)(17), P(5)(19), P(4)(21), Sum(92), Cout(92));
FA74 : full_adder port map(P(3)(23), P(2)(25), P(1)(27), Sum(93), Cout(93));
FA75 : full_adder port map(P(0)(29), Cout(6), Cout(7), Sum(94), Cout(94));
FA76 : full_adder port map(Cout(8), Sum(9), Sum(10), Sum(95), Cout(95));
FA77 : full_adder port map(P(5)(20), P(4)(22), P(3)(24), Sum(96), Cout(96));
FA78 : full_adder port map(P(2)(26), P(1)(28), P(0)(30), Sum(97), Cout(97));
FA79 : full_adder port map(Cout(9), Cout(10), Cout(11), Sum(98), Cout(98));
FA80 : full_adder port map(Sum(12), Sum(13), Sum(14), Sum(99), Cout(99));
FA81 : full_adder port map(P(4)(23), P(3)(25), P(2)(27), Sum(100), Cout(100));
FA82 : full_adder port map(P(1)(29), P(0)(31), Cout(12), Sum(101), Cout(101));
FA83 : full_adder port map(Cout(13), Cout(14), Cout(15), Sum(102), Cout(102));
FA84 : full_adder port map(Sum(16), Sum(17), Sum(18), Sum(103), Cout(103));
FA85 : full_adder port map(P(4)(24), P(3)(26), P(2)(28), Sum(104), Cout(104));
FA86 : full_adder port map(P(1)(30), P(0)(32), Cout(16), Sum(105), Cout(105));
FA87 : full_adder port map(Cout(17), Cout(18), Cout(19), Sum(106), Cout(106));
FA88 : full_adder port map(Sum(20), Sum(21), Sum(22), Sum(107), Cout(107));
FA89 : full_adder port map(P(12)(9), P(13)(7), P(14)(5), Sum(108), Cout(108));
FA90 : full_adder port map(P(15)(3), P(16)(1), Cout(20), Sum(109), Cout(109));
FA91 : full_adder port map(Cout(21), Cout(22), Cout(23), Sum(110), Cout(110));
FA92 : full_adder port map(Sum(24), Sum(25), Sum(26), Sum(111), Cout(111));
FA93 : full_adder port map(P(12)(10), P(13)(8), P(14)(6), Sum(112), Cout(112));
FA94 : full_adder port map(P(15)(4), P(16)(2), Cout(24), Sum(113), Cout(113));
FA95 : full_adder port map(Cout(25), Cout(26), Cout(27), Sum(114), Cout(114));
FA96 : full_adder port map(Sum(28), Sum(29), Sum(30), Sum(115), Cout(115));
FA97 : full_adder port map(P(12)(11), P(13)(9), P(14)(7), Sum(116), Cout(116));
FA98 : full_adder port map(P(15)(5), P(16)(3), Cout(28), Sum(117), Cout(117));
FA99 : full_adder port map(Cout(29), Cout(30), Cout(31), Sum(118), Cout(118));
FA100 : full_adder port map(Sum(32), Sum(33), Sum(34), Sum(119), Cout(119));
FA101 : full_adder port map(P(12)(12), P(13)(10), P(14)(8), Sum(120), Cout(120));
FA102 : full_adder port map(P(15)(6), P(16)(4), Cout(32), Sum(121), Cout(121));
FA103 : full_adder port map(Cout(33), Cout(34), Cout(35), Sum(122), Cout(122));
FA104 : full_adder port map(Sum(36), Sum(37), Sum(38), Sum(123), Cout(123));
FA105 : full_adder port map(P(11)(15), P(12)(13), P(13)(11), Sum(124), Cout(124));
FA106 : full_adder port map(P(14)(9), P(15)(7), P(16)(5), Sum(125), Cout(125));
FA107 : full_adder port map(Cout(36), Cout(37), Cout(38), Sum(126), Cout(126));
FA108 : full_adder port map(Cout(39), Sum(40), Sum(41), Sum(127), Cout(127));
FA109 : full_adder port map(P(10)(18), P(11)(16), P(12)(14), Sum(128), Cout(128));
FA110 : full_adder port map(P(13)(12), P(14)(10), P(15)(8), Sum(129), Cout(129));
FA111 : full_adder port map(P(16)(6), Cout(40), Cout(41), Sum(130), Cout(130));
FA112 : full_adder port map(Cout(42), Sum(43), Sum(44), Sum(131), Cout(131));
FA113 : full_adder port map(P(9)(21), P(10)(19), P(11)(17), Sum(132), Cout(132));
FA114 : full_adder port map(P(12)(15), P(13)(13), P(14)(11), Sum(133), Cout(133));
FA115 : full_adder port map(P(15)(9), P(16)(7), Cout(43), Sum(134), Cout(134));
FA116 : full_adder port map(Cout(44), Cout(45), Sum(46), Sum(135), Cout(135));
FA117 : full_adder port map(P(8)(24), P(9)(22), P(10)(20), Sum(136), Cout(136));
FA118 : full_adder port map(P(11)(18), P(12)(16), P(13)(14), Sum(137), Cout(137));
FA119 : full_adder port map(P(14)(12), P(15)(10), P(16)(8), Sum(138), Cout(138));
FA120 : full_adder port map(Cout(46), Cout(47), Sum(48), Sum(139), Cout(139));
FA121 : full_adder port map(P(7)(27), P(8)(25), P(9)(23), Sum(140), Cout(140));
FA122 : full_adder port map(P(10)(21), P(11)(19), P(12)(17), Sum(141), Cout(141));
FA123 : full_adder port map(P(13)(15), P(14)(13), P(15)(11), Sum(142), Cout(142));
FA124 : full_adder port map(P(16)(9), Cout(48), Cout(49), Sum(143), Cout(143));
FA125 : full_adder port map(P(6)(30), P(7)(28), P(8)(26), Sum(144), Cout(144));
FA126 : full_adder port map(P(9)(24), P(10)(22), P(11)(20), Sum(145), Cout(145));
FA127 : full_adder port map(P(12)(18), P(13)(16), P(14)(14), Sum(146), Cout(146));
FA128 : full_adder port map(P(15)(12), P(16)(10), Cout(50), Sum(147), Cout(147));
FA129 : full_adder port map(nSig(5), P(6)(31), P(7)(29), Sum(148), Cout(148));
FA130 : full_adder port map(P(8)(27), P(9)(25), P(10)(23), Sum(149), Cout(149));
FA131 : full_adder port map(P(11)(21), P(12)(19), P(13)(17), Sum(150), Cout(150));
FA132 : full_adder port map(P(14)(15), P(15)(13), P(16)(11), Sum(151), Cout(151));
FA133 : full_adder port map('1', P(6)(32), P(7)(30), Sum(152), Cout(152));
FA134 : full_adder port map(P(8)(28), P(9)(26), P(10)(24), Sum(153), Cout(153));
FA135 : full_adder port map(P(11)(22), P(12)(20), P(13)(18), Sum(154), Cout(154));
HA21 : half_adder port map(P(14)(16), P(15)(14), Sum(155), Cout(155));
FA136 : full_adder port map(nSig(6), P(7)(31), P(8)(29), Sum(156), Cout(156));
FA137 : full_adder port map(P(9)(27), P(10)(25), P(11)(23), Sum(157), Cout(157));
FA138 : full_adder port map(P(12)(21), P(13)(19), P(14)(17), Sum(158), Cout(158));
FA139 : full_adder port map('1', P(7)(32), P(8)(30), Sum(159), Cout(159));
FA140 : full_adder port map(P(9)(28), P(10)(26), P(11)(24), Sum(160), Cout(160));
HA22 : half_adder port map(P(12)(22), P(13)(20), Sum(161), Cout(161));
FA141 : full_adder port map(nSig(7), P(8)(31), P(9)(29), Sum(162), Cout(162));
FA142 : full_adder port map(P(10)(27), P(11)(25), P(12)(23), Sum(163), Cout(163));
FA143 : full_adder port map('1', P(8)(32), P(9)(30), Sum(164), Cout(164));
HA23 : half_adder port map(P(10)(28), P(11)(26), Sum(165), Cout(165));
FA144 : full_adder port map(nSig(8), P(9)(31), P(10)(29), Sum(166), Cout(166));
HA24 : half_adder port map('1', P(9)(32), Sum(167), Cout(167));
HA25 : half_adder port map(Sig(5), P(5)(0), Sum(168), Cout(168));
HA26 : half_adder port map(P(5)(1), P(4)(3), Sum(169), Cout(169));
FA145 : full_adder port map(Sig(6), P(6)(0), P(5)(2), Sum(170), Cout(170));
HA27 : half_adder port map(P(4)(4), P(3)(6), Sum(171), Cout(171));
FA146 : full_adder port map(P(6)(1), P(5)(3), P(4)(5), Sum(172), Cout(172));
HA28 : half_adder port map(P(3)(7), P(2)(9), Sum(173), Cout(173));
FA147 : full_adder port map(Sig(7), P(7)(0), P(6)(2), Sum(174), Cout(174));
FA148 : full_adder port map(P(5)(4), P(4)(6), P(3)(8), Sum(175), Cout(175));
HA29 : half_adder port map(P(2)(10), P(1)(12), Sum(176), Cout(176));
FA149 : full_adder port map(P(7)(1), P(6)(3), P(5)(5), Sum(177), Cout(177));
FA150 : full_adder port map(P(4)(7), P(3)(9), P(2)(11), Sum(178), Cout(178));
HA30 : half_adder port map(P(1)(13), P(0)(15), Sum(179), Cout(179));
FA151 : full_adder port map(P(7)(2), P(6)(4), P(5)(6), Sum(180), Cout(180));
FA152 : full_adder port map(P(4)(8), P(3)(10), P(2)(12), Sum(181), Cout(181));
FA153 : full_adder port map(P(1)(14), P(0)(16), Sum(52), Sum(182), Cout(182));
FA154 : full_adder port map(P(6)(5), P(5)(7), P(4)(9), Sum(183), Cout(183));
FA155 : full_adder port map(P(3)(11), P(2)(13), P(1)(15), Sum(184), Cout(184));
FA156 : full_adder port map(P(0)(17), Cout(52), Sum(53), Sum(185), Cout(185));
FA157 : full_adder port map(P(5)(8), P(4)(10), P(3)(12), Sum(186), Cout(186));
FA158 : full_adder port map(P(2)(14), P(1)(16), P(0)(18), Sum(187), Cout(187));
FA159 : full_adder port map(Cout(53), Sum(54), Sum(55), Sum(188), Cout(188));
FA160 : full_adder port map(P(4)(11), P(3)(13), P(2)(15), Sum(189), Cout(189));
FA161 : full_adder port map(P(1)(17), P(0)(19), Cout(54), Sum(190), Cout(190));
FA162 : full_adder port map(Cout(55), Sum(56), Sum(57), Sum(191), Cout(191));
FA163 : full_adder port map(P(3)(14), P(2)(16), P(1)(18), Sum(192), Cout(192));
FA164 : full_adder port map(P(0)(20), Cout(56), Cout(57), Sum(193), Cout(193));
FA165 : full_adder port map(Sum(58), Sum(59), Sum(60), Sum(194), Cout(194));
FA166 : full_adder port map(P(2)(17), P(1)(19), P(0)(21), Sum(195), Cout(195));
FA167 : full_adder port map(Cout(58), Cout(59), Cout(60), Sum(196), Cout(196));
FA168 : full_adder port map(Sum(61), Sum(62), Sum(63), Sum(197), Cout(197));
FA169 : full_adder port map(P(1)(20), P(0)(22), Cout(61), Sum(198), Cout(198));
FA170 : full_adder port map(Cout(62), Cout(63), Sum(64), Sum(199), Cout(199));
FA171 : full_adder port map(Sum(65), Sum(66), Sum(67), Sum(200), Cout(200));
FA172 : full_adder port map(P(0)(23), Cout(64), Cout(65), Sum(201), Cout(201));
FA173 : full_adder port map(Cout(66), Cout(67), Sum(68), Sum(202), Cout(202));
FA174 : full_adder port map(Sum(69), Sum(70), Sum(71), Sum(203), Cout(203));
FA175 : full_adder port map(Sum(0), Cout(68), Cout(69), Sum(204), Cout(204));
FA176 : full_adder port map(Cout(70), Cout(71), Sum(72), Sum(205), Cout(205));
FA177 : full_adder port map(Sum(73), Sum(74), Sum(75), Sum(206), Cout(206));
FA178 : full_adder port map(Sum(1), Cout(72), Cout(73), Sum(207), Cout(207));
FA179 : full_adder port map(Cout(74), Cout(75), Sum(76), Sum(208), Cout(208));
FA180 : full_adder port map(Sum(77), Sum(78), Sum(79), Sum(209), Cout(209));
FA181 : full_adder port map(Sum(3), Cout(76), Cout(77), Sum(210), Cout(210));
FA182 : full_adder port map(Cout(78), Cout(79), Sum(80), Sum(211), Cout(211));
FA183 : full_adder port map(Sum(81), Sum(82), Sum(83), Sum(212), Cout(212));
FA184 : full_adder port map(Sum(5), Cout(80), Cout(81), Sum(213), Cout(213));
FA185 : full_adder port map(Cout(82), Cout(83), Sum(84), Sum(214), Cout(214));
FA186 : full_adder port map(Sum(85), Sum(86), Sum(87), Sum(215), Cout(215));
FA187 : full_adder port map(Sum(8), Cout(84), Cout(85), Sum(216), Cout(216));
FA188 : full_adder port map(Cout(86), Cout(87), Sum(88), Sum(217), Cout(217));
FA189 : full_adder port map(Sum(89), Sum(90), Sum(91), Sum(218), Cout(218));
FA190 : full_adder port map(Sum(11), Cout(88), Cout(89), Sum(219), Cout(219));
FA191 : full_adder port map(Cout(90), Cout(91), Sum(92), Sum(220), Cout(220));
FA192 : full_adder port map(Sum(93), Sum(94), Sum(95), Sum(221), Cout(221));
FA193 : full_adder port map(Sum(15), Cout(92), Cout(93), Sum(222), Cout(222));
FA194 : full_adder port map(Cout(94), Cout(95), Sum(96), Sum(223), Cout(223));
FA195 : full_adder port map(Sum(97), Sum(98), Sum(99), Sum(224), Cout(224));
FA196 : full_adder port map(Sum(19), Cout(96), Cout(97), Sum(225), Cout(225));
FA197 : full_adder port map(Cout(98), Cout(99), Sum(100), Sum(226), Cout(226));
FA198 : full_adder port map(Sum(101), Sum(102), Sum(103), Sum(227), Cout(227));
FA199 : full_adder port map(Sum(23), Cout(100), Cout(101), Sum(228), Cout(228));
FA200 : full_adder port map(Cout(102), Cout(103), Sum(104), Sum(229), Cout(229));
FA201 : full_adder port map(Sum(105), Sum(106), Sum(107), Sum(230), Cout(230));
FA202 : full_adder port map(Sum(27), Cout(104), Cout(105), Sum(231), Cout(231));
FA203 : full_adder port map(Cout(106), Cout(107), Sum(108), Sum(232), Cout(232));
FA204 : full_adder port map(Sum(109), Sum(110), Sum(111), Sum(233), Cout(233));
FA205 : full_adder port map(Sum(31), Cout(108), Cout(109), Sum(234), Cout(234));
FA206 : full_adder port map(Cout(110), Cout(111), Sum(112), Sum(235), Cout(235));
FA207 : full_adder port map(Sum(113), Sum(114), Sum(115), Sum(236), Cout(236));
FA208 : full_adder port map(Sum(35), Cout(112), Cout(113), Sum(237), Cout(237));
FA209 : full_adder port map(Cout(114), Cout(115), Sum(116), Sum(238), Cout(238));
FA210 : full_adder port map(Sum(117), Sum(118), Sum(119), Sum(239), Cout(239));
FA211 : full_adder port map(Sum(39), Cout(116), Cout(117), Sum(240), Cout(240));
FA212 : full_adder port map(Cout(118), Cout(119), Sum(120), Sum(241), Cout(241));
FA213 : full_adder port map(Sum(121), Sum(122), Sum(123), Sum(242), Cout(242));
FA214 : full_adder port map(Sum(42), Cout(120), Cout(121), Sum(243), Cout(243));
FA215 : full_adder port map(Cout(122), Cout(123), Sum(124), Sum(244), Cout(244));
FA216 : full_adder port map(Sum(125), Sum(126), Sum(127), Sum(245), Cout(245));
FA217 : full_adder port map(Sum(45), Cout(124), Cout(125), Sum(246), Cout(246));
FA218 : full_adder port map(Cout(126), Cout(127), Sum(128), Sum(247), Cout(247));
FA219 : full_adder port map(Sum(129), Sum(130), Sum(131), Sum(248), Cout(248));
FA220 : full_adder port map(Sum(47), Cout(128), Cout(129), Sum(249), Cout(249));
FA221 : full_adder port map(Cout(130), Cout(131), Sum(132), Sum(250), Cout(250));
FA222 : full_adder port map(Sum(133), Sum(134), Sum(135), Sum(251), Cout(251));
FA223 : full_adder port map(Sum(49), Cout(132), Cout(133), Sum(252), Cout(252));
FA224 : full_adder port map(Cout(134), Cout(135), Sum(136), Sum(253), Cout(253));
FA225 : full_adder port map(Sum(137), Sum(138), Sum(139), Sum(254), Cout(254));
FA226 : full_adder port map(Sum(50), Cout(136), Cout(137), Sum(255), Cout(255));
FA227 : full_adder port map(Cout(138), Cout(139), Sum(140), Sum(256), Cout(256));
FA228 : full_adder port map(Sum(141), Sum(142), Sum(143), Sum(257), Cout(257));
FA229 : full_adder port map(Sum(51), Cout(140), Cout(141), Sum(258), Cout(258));
FA230 : full_adder port map(Cout(142), Cout(143), Sum(144), Sum(259), Cout(259));
FA231 : full_adder port map(Sum(145), Sum(146), Sum(147), Sum(260), Cout(260));
FA232 : full_adder port map(Cout(51), Cout(144), Cout(145), Sum(261), Cout(261));
FA233 : full_adder port map(Cout(146), Cout(147), Sum(148), Sum(262), Cout(262));
FA234 : full_adder port map(Sum(149), Sum(150), Sum(151), Sum(263), Cout(263));
FA235 : full_adder port map(P(16)(12), Cout(148), Cout(149), Sum(264), Cout(264));
FA236 : full_adder port map(Cout(150), Cout(151), Sum(152), Sum(265), Cout(265));
FA237 : full_adder port map(Sum(153), Sum(154), Sum(155), Sum(266), Cout(266));
FA238 : full_adder port map(P(15)(15), P(16)(13), Cout(152), Sum(267), Cout(267));
FA239 : full_adder port map(Cout(153), Cout(154), Cout(155), Sum(268), Cout(268));
FA240 : full_adder port map(Sum(156), Sum(157), Sum(158), Sum(269), Cout(269));
FA241 : full_adder port map(P(14)(18), P(15)(16), P(16)(14), Sum(270), Cout(270));
FA242 : full_adder port map(Cout(156), Cout(157), Cout(158), Sum(271), Cout(271));
FA243 : full_adder port map(Sum(159), Sum(160), Sum(161), Sum(272), Cout(272));
FA244 : full_adder port map(P(13)(21), P(14)(19), P(15)(17), Sum(273), Cout(273));
FA245 : full_adder port map(P(16)(15), Cout(159), Cout(160), Sum(274), Cout(274));
FA246 : full_adder port map(Cout(161), Sum(162), Sum(163), Sum(275), Cout(275));
FA247 : full_adder port map(P(12)(24), P(13)(22), P(14)(20), Sum(276), Cout(276));
FA248 : full_adder port map(P(15)(18), P(16)(16), Cout(162), Sum(277), Cout(277));
FA249 : full_adder port map(Cout(163), Sum(164), Sum(165), Sum(278), Cout(278));
FA250 : full_adder port map(P(11)(27), P(12)(25), P(13)(23), Sum(279), Cout(279));
FA251 : full_adder port map(P(14)(21), P(15)(19), P(16)(17), Sum(280), Cout(280));
FA252 : full_adder port map(Cout(164), Cout(165), Sum(166), Sum(281), Cout(281));
FA253 : full_adder port map(P(10)(30), P(11)(28), P(12)(26), Sum(282), Cout(282));
FA254 : full_adder port map(P(13)(24), P(14)(22), P(15)(20), Sum(283), Cout(283));
FA255 : full_adder port map(P(16)(18), Cout(166), Sum(167), Sum(284), Cout(284));
FA256 : full_adder port map(nSig(9), P(10)(31), P(11)(29), Sum(285), Cout(285));
FA257 : full_adder port map(P(12)(27), P(13)(25), P(14)(23), Sum(286), Cout(286));
FA258 : full_adder port map(P(15)(21), P(16)(19), Cout(167), Sum(287), Cout(287));
FA259 : full_adder port map('1', P(10)(32), P(11)(30), Sum(288), Cout(288));
FA260 : full_adder port map(P(12)(28), P(13)(26), P(14)(24), Sum(289), Cout(289));
HA31 : half_adder port map(P(15)(22), P(16)(20), Sum(290), Cout(290));
FA261 : full_adder port map(nSig(10), P(11)(31), P(12)(29), Sum(291), Cout(291));
FA262 : full_adder port map(P(13)(27), P(14)(25), P(15)(23), Sum(292), Cout(292));
FA263 : full_adder port map('1', P(11)(32), P(12)(30), Sum(293), Cout(293));
HA32 : half_adder port map(P(13)(28), P(14)(26), Sum(294), Cout(294));
FA264 : full_adder port map(nSig(11), P(12)(31), P(13)(29), Sum(295), Cout(295));
HA33 : half_adder port map('1', P(12)(32), Sum(296), Cout(296));
HA34 : half_adder port map(Sig(3), P(3)(0), Sum(297), Cout(297));
HA35 : half_adder port map(P(3)(1), P(2)(3), Sum(298), Cout(298));
FA265 : full_adder port map(Sig(4), P(4)(0), P(3)(2), Sum(299), Cout(299));
HA36 : half_adder port map(P(2)(4), P(1)(6), Sum(300), Cout(300));
FA266 : full_adder port map(P(4)(1), P(3)(3), P(2)(5), Sum(301), Cout(301));
HA37 : half_adder port map(P(1)(7), P(0)(9), Sum(302), Cout(302));
FA267 : full_adder port map(P(4)(2), P(3)(4), P(2)(6), Sum(303), Cout(303));
FA268 : full_adder port map(P(1)(8), P(0)(10), Sum(168), Sum(304), Cout(304));
FA269 : full_adder port map(P(3)(5), P(2)(7), P(1)(9), Sum(305), Cout(305));
FA270 : full_adder port map(P(0)(11), Cout(168), Sum(169), Sum(306), Cout(306));
FA271 : full_adder port map(P(2)(8), P(1)(10), P(0)(12), Sum(307), Cout(307));
FA272 : full_adder port map(Cout(169), Sum(170), Sum(171), Sum(308), Cout(308));
FA273 : full_adder port map(P(1)(11), P(0)(13), Cout(170), Sum(309), Cout(309));
FA274 : full_adder port map(Cout(171), Sum(172), Sum(173), Sum(310), Cout(310));
FA275 : full_adder port map(P(0)(14), Cout(172), Cout(173), Sum(311), Cout(311));
FA276 : full_adder port map(Sum(174), Sum(175), Sum(176), Sum(312), Cout(312));
FA277 : full_adder port map(Cout(174), Cout(175), Cout(176), Sum(313), Cout(313));
FA278 : full_adder port map(Sum(177), Sum(178), Sum(179), Sum(314), Cout(314));
FA279 : full_adder port map(Cout(177), Cout(178), Cout(179), Sum(315), Cout(315));
FA280 : full_adder port map(Sum(180), Sum(181), Sum(182), Sum(316), Cout(316));
FA281 : full_adder port map(Cout(180), Cout(181), Cout(182), Sum(317), Cout(317));
FA282 : full_adder port map(Sum(183), Sum(184), Sum(185), Sum(318), Cout(318));
FA283 : full_adder port map(Cout(183), Cout(184), Cout(185), Sum(319), Cout(319));
FA284 : full_adder port map(Sum(186), Sum(187), Sum(188), Sum(320), Cout(320));
FA285 : full_adder port map(Cout(186), Cout(187), Cout(188), Sum(321), Cout(321));
FA286 : full_adder port map(Sum(189), Sum(190), Sum(191), Sum(322), Cout(322));
FA287 : full_adder port map(Cout(189), Cout(190), Cout(191), Sum(323), Cout(323));
FA288 : full_adder port map(Sum(192), Sum(193), Sum(194), Sum(324), Cout(324));
FA289 : full_adder port map(Cout(192), Cout(193), Cout(194), Sum(325), Cout(325));
FA290 : full_adder port map(Sum(195), Sum(196), Sum(197), Sum(326), Cout(326));
FA291 : full_adder port map(Cout(195), Cout(196), Cout(197), Sum(327), Cout(327));
FA292 : full_adder port map(Sum(198), Sum(199), Sum(200), Sum(328), Cout(328));
FA293 : full_adder port map(Cout(198), Cout(199), Cout(200), Sum(329), Cout(329));
FA294 : full_adder port map(Sum(201), Sum(202), Sum(203), Sum(330), Cout(330));
FA295 : full_adder port map(Cout(201), Cout(202), Cout(203), Sum(331), Cout(331));
FA296 : full_adder port map(Sum(204), Sum(205), Sum(206), Sum(332), Cout(332));
FA297 : full_adder port map(Cout(204), Cout(205), Cout(206), Sum(333), Cout(333));
FA298 : full_adder port map(Sum(207), Sum(208), Sum(209), Sum(334), Cout(334));
FA299 : full_adder port map(Cout(207), Cout(208), Cout(209), Sum(335), Cout(335));
FA300 : full_adder port map(Sum(210), Sum(211), Sum(212), Sum(336), Cout(336));
FA301 : full_adder port map(Cout(210), Cout(211), Cout(212), Sum(337), Cout(337));
FA302 : full_adder port map(Sum(213), Sum(214), Sum(215), Sum(338), Cout(338));
FA303 : full_adder port map(Cout(213), Cout(214), Cout(215), Sum(339), Cout(339));
FA304 : full_adder port map(Sum(216), Sum(217), Sum(218), Sum(340), Cout(340));
FA305 : full_adder port map(Cout(216), Cout(217), Cout(218), Sum(341), Cout(341));
FA306 : full_adder port map(Sum(219), Sum(220), Sum(221), Sum(342), Cout(342));
FA307 : full_adder port map(Cout(219), Cout(220), Cout(221), Sum(343), Cout(343));
FA308 : full_adder port map(Sum(222), Sum(223), Sum(224), Sum(344), Cout(344));
FA309 : full_adder port map(Cout(222), Cout(223), Cout(224), Sum(345), Cout(345));
FA310 : full_adder port map(Sum(225), Sum(226), Sum(227), Sum(346), Cout(346));
FA311 : full_adder port map(Cout(225), Cout(226), Cout(227), Sum(347), Cout(347));
FA312 : full_adder port map(Sum(228), Sum(229), Sum(230), Sum(348), Cout(348));
FA313 : full_adder port map(Cout(228), Cout(229), Cout(230), Sum(349), Cout(349));
FA314 : full_adder port map(Sum(231), Sum(232), Sum(233), Sum(350), Cout(350));
FA315 : full_adder port map(Cout(231), Cout(232), Cout(233), Sum(351), Cout(351));
FA316 : full_adder port map(Sum(234), Sum(235), Sum(236), Sum(352), Cout(352));
FA317 : full_adder port map(Cout(234), Cout(235), Cout(236), Sum(353), Cout(353));
FA318 : full_adder port map(Sum(237), Sum(238), Sum(239), Sum(354), Cout(354));
FA319 : full_adder port map(Cout(237), Cout(238), Cout(239), Sum(355), Cout(355));
FA320 : full_adder port map(Sum(240), Sum(241), Sum(242), Sum(356), Cout(356));
FA321 : full_adder port map(Cout(240), Cout(241), Cout(242), Sum(357), Cout(357));
FA322 : full_adder port map(Sum(243), Sum(244), Sum(245), Sum(358), Cout(358));
FA323 : full_adder port map(Cout(243), Cout(244), Cout(245), Sum(359), Cout(359));
FA324 : full_adder port map(Sum(246), Sum(247), Sum(248), Sum(360), Cout(360));
FA325 : full_adder port map(Cout(246), Cout(247), Cout(248), Sum(361), Cout(361));
FA326 : full_adder port map(Sum(249), Sum(250), Sum(251), Sum(362), Cout(362));
FA327 : full_adder port map(Cout(249), Cout(250), Cout(251), Sum(363), Cout(363));
FA328 : full_adder port map(Sum(252), Sum(253), Sum(254), Sum(364), Cout(364));
FA329 : full_adder port map(Cout(252), Cout(253), Cout(254), Sum(365), Cout(365));
FA330 : full_adder port map(Sum(255), Sum(256), Sum(257), Sum(366), Cout(366));
FA331 : full_adder port map(Cout(255), Cout(256), Cout(257), Sum(367), Cout(367));
FA332 : full_adder port map(Sum(258), Sum(259), Sum(260), Sum(368), Cout(368));
FA333 : full_adder port map(Cout(258), Cout(259), Cout(260), Sum(369), Cout(369));
FA334 : full_adder port map(Sum(261), Sum(262), Sum(263), Sum(370), Cout(370));
FA335 : full_adder port map(Cout(261), Cout(262), Cout(263), Sum(371), Cout(371));
FA336 : full_adder port map(Sum(264), Sum(265), Sum(266), Sum(372), Cout(372));
FA337 : full_adder port map(Cout(264), Cout(265), Cout(266), Sum(373), Cout(373));
FA338 : full_adder port map(Sum(267), Sum(268), Sum(269), Sum(374), Cout(374));
FA339 : full_adder port map(Cout(267), Cout(268), Cout(269), Sum(375), Cout(375));
FA340 : full_adder port map(Sum(270), Sum(271), Sum(272), Sum(376), Cout(376));
FA341 : full_adder port map(Cout(270), Cout(271), Cout(272), Sum(377), Cout(377));
FA342 : full_adder port map(Sum(273), Sum(274), Sum(275), Sum(378), Cout(378));
FA343 : full_adder port map(Cout(273), Cout(274), Cout(275), Sum(379), Cout(379));
FA344 : full_adder port map(Sum(276), Sum(277), Sum(278), Sum(380), Cout(380));
FA345 : full_adder port map(Cout(276), Cout(277), Cout(278), Sum(381), Cout(381));
FA346 : full_adder port map(Sum(279), Sum(280), Sum(281), Sum(382), Cout(382));
FA347 : full_adder port map(Cout(279), Cout(280), Cout(281), Sum(383), Cout(383));
FA348 : full_adder port map(Sum(282), Sum(283), Sum(284), Sum(384), Cout(384));
FA349 : full_adder port map(Cout(282), Cout(283), Cout(284), Sum(385), Cout(385));
FA350 : full_adder port map(Sum(285), Sum(286), Sum(287), Sum(386), Cout(386));
FA351 : full_adder port map(Cout(285), Cout(286), Cout(287), Sum(387), Cout(387));
FA352 : full_adder port map(Sum(288), Sum(289), Sum(290), Sum(388), Cout(388));
FA353 : full_adder port map(P(16)(21), Cout(288), Cout(289), Sum(389), Cout(389));
FA354 : full_adder port map(Cout(290), Sum(291), Sum(292), Sum(390), Cout(390));
FA355 : full_adder port map(P(15)(24), P(16)(22), Cout(291), Sum(391), Cout(391));
FA356 : full_adder port map(Cout(292), Sum(293), Sum(294), Sum(392), Cout(392));
FA357 : full_adder port map(P(14)(27), P(15)(25), P(16)(23), Sum(393), Cout(393));
FA358 : full_adder port map(Cout(293), Cout(294), Sum(295), Sum(394), Cout(394));
FA359 : full_adder port map(P(13)(30), P(14)(28), P(15)(26), Sum(395), Cout(395));
FA360 : full_adder port map(P(16)(24), Cout(295), Sum(296), Sum(396), Cout(396));
FA361 : full_adder port map(nSig(12), P(13)(31), P(14)(29), Sum(397), Cout(397));
FA362 : full_adder port map(P(15)(27), P(16)(25), Cout(296), Sum(398), Cout(398));
FA363 : full_adder port map('1', P(13)(32), P(14)(30), Sum(399), Cout(399));
HA38 : half_adder port map(P(15)(28), P(16)(26), Sum(400), Cout(400));
FA364 : full_adder port map(nSig(13), P(14)(31), P(15)(29), Sum(401), Cout(401));
HA39 : half_adder port map('1', P(14)(32), Sum(402), Cout(402));
HA40 : half_adder port map(Sig(2), P(2)(0), Sum(403), Cout(403));
HA41 : half_adder port map(P(2)(1), P(1)(3), Sum(404), Cout(404));
FA365 : full_adder port map(P(2)(2), P(1)(4), P(0)(6), Sum(405), Cout(405));
FA366 : full_adder port map(P(1)(5), P(0)(7), Cout(297), Sum(406), Cout(406));
FA367 : full_adder port map(P(0)(8), Cout(298), Sum(299), Sum(407), Cout(407));
FA368 : full_adder port map(Cout(299), Cout(300), Sum(301), Sum(408), Cout(408));
FA369 : full_adder port map(Cout(301), Cout(302), Sum(303), Sum(409), Cout(409));
FA370 : full_adder port map(Cout(303), Cout(304), Sum(305), Sum(410), Cout(410));
FA371 : full_adder port map(Cout(305), Cout(306), Sum(307), Sum(411), Cout(411));
FA372 : full_adder port map(Cout(307), Cout(308), Sum(309), Sum(412), Cout(412));
FA373 : full_adder port map(Cout(309), Cout(310), Sum(311), Sum(413), Cout(413));
FA374 : full_adder port map(Cout(311), Cout(312), Sum(313), Sum(414), Cout(414));
FA375 : full_adder port map(Cout(313), Cout(314), Sum(315), Sum(415), Cout(415));
FA376 : full_adder port map(Cout(315), Cout(316), Sum(317), Sum(416), Cout(416));
FA377 : full_adder port map(Cout(317), Cout(318), Sum(319), Sum(417), Cout(417));
FA378 : full_adder port map(Cout(319), Cout(320), Sum(321), Sum(418), Cout(418));
FA379 : full_adder port map(Cout(321), Cout(322), Sum(323), Sum(419), Cout(419));
FA380 : full_adder port map(Cout(323), Cout(324), Sum(325), Sum(420), Cout(420));
FA381 : full_adder port map(Cout(325), Cout(326), Sum(327), Sum(421), Cout(421));
FA382 : full_adder port map(Cout(327), Cout(328), Sum(329), Sum(422), Cout(422));
FA383 : full_adder port map(Cout(329), Cout(330), Sum(331), Sum(423), Cout(423));
FA384 : full_adder port map(Cout(331), Cout(332), Sum(333), Sum(424), Cout(424));
FA385 : full_adder port map(Cout(333), Cout(334), Sum(335), Sum(425), Cout(425));
FA386 : full_adder port map(Cout(335), Cout(336), Sum(337), Sum(426), Cout(426));
FA387 : full_adder port map(Cout(337), Cout(338), Sum(339), Sum(427), Cout(427));
FA388 : full_adder port map(Cout(339), Cout(340), Sum(341), Sum(428), Cout(428));
FA389 : full_adder port map(Cout(341), Cout(342), Sum(343), Sum(429), Cout(429));
FA390 : full_adder port map(Cout(343), Cout(344), Sum(345), Sum(430), Cout(430));
FA391 : full_adder port map(Cout(345), Cout(346), Sum(347), Sum(431), Cout(431));
FA392 : full_adder port map(Cout(347), Cout(348), Sum(349), Sum(432), Cout(432));
FA393 : full_adder port map(Cout(349), Cout(350), Sum(351), Sum(433), Cout(433));
FA394 : full_adder port map(Cout(351), Cout(352), Sum(353), Sum(434), Cout(434));
FA395 : full_adder port map(Cout(353), Cout(354), Sum(355), Sum(435), Cout(435));
FA396 : full_adder port map(Cout(355), Cout(356), Sum(357), Sum(436), Cout(436));
FA397 : full_adder port map(Cout(357), Cout(358), Sum(359), Sum(437), Cout(437));
FA398 : full_adder port map(Cout(359), Cout(360), Sum(361), Sum(438), Cout(438));
FA399 : full_adder port map(Cout(361), Cout(362), Sum(363), Sum(439), Cout(439));
FA400 : full_adder port map(Cout(363), Cout(364), Sum(365), Sum(440), Cout(440));
FA401 : full_adder port map(Cout(365), Cout(366), Sum(367), Sum(441), Cout(441));
FA402 : full_adder port map(Cout(367), Cout(368), Sum(369), Sum(442), Cout(442));
FA403 : full_adder port map(Cout(369), Cout(370), Sum(371), Sum(443), Cout(443));
FA404 : full_adder port map(Cout(371), Cout(372), Sum(373), Sum(444), Cout(444));
FA405 : full_adder port map(Cout(373), Cout(374), Sum(375), Sum(445), Cout(445));
FA406 : full_adder port map(Cout(375), Cout(376), Sum(377), Sum(446), Cout(446));
FA407 : full_adder port map(Cout(377), Cout(378), Sum(379), Sum(447), Cout(447));
FA408 : full_adder port map(Cout(379), Cout(380), Sum(381), Sum(448), Cout(448));
FA409 : full_adder port map(Cout(381), Cout(382), Sum(383), Sum(449), Cout(449));
FA410 : full_adder port map(Cout(383), Cout(384), Sum(385), Sum(450), Cout(450));
FA411 : full_adder port map(Cout(385), Cout(386), Sum(387), Sum(451), Cout(451));
FA412 : full_adder port map(Cout(387), Cout(388), Sum(389), Sum(452), Cout(452));
FA413 : full_adder port map(Cout(389), Cout(390), Sum(391), Sum(453), Cout(453));
FA414 : full_adder port map(Cout(391), Cout(392), Sum(393), Sum(454), Cout(454));
FA415 : full_adder port map(Cout(393), Cout(394), Sum(395), Sum(455), Cout(455));
FA416 : full_adder port map(Cout(395), Cout(396), Sum(397), Sum(456), Cout(456));
FA417 : full_adder port map(Cout(397), Cout(398), Sum(399), Sum(457), Cout(457));
FA418 : full_adder port map(P(16)(27), Cout(399), Cout(400), Sum(458), Cout(458));
FA419 : full_adder port map(P(15)(30), P(16)(28), Cout(401), Sum(459), Cout(459));
FA420 : full_adder port map(nSig(14), P(15)(31), P(16)(29), Sum(460), Cout(460));
HA42 : half_adder port map('1', P(15)(32), Sum(461), Cout(461));
HA43 : half_adder port map(Sig(1), P(1)(0), Sum(462), Cout(462));
HA44 : half_adder port map(P(1)(1), P(0)(3), Sum(463), Cout(463));
FA421 : full_adder port map(P(1)(2), P(0)(4), Sum(403), Sum(464), Cout(464));
FA422 : full_adder port map(P(0)(5), Cout(403), Sum(404), Sum(465), Cout(465));
FA423 : full_adder port map(Sum(297), Cout(404), Sum(405), Sum(466), Cout(466));
FA424 : full_adder port map(Sum(298), Cout(405), Sum(406), Sum(467), Cout(467));
FA425 : full_adder port map(Sum(300), Cout(406), Sum(407), Sum(468), Cout(468));
FA426 : full_adder port map(Sum(302), Cout(407), Sum(408), Sum(469), Cout(469));
FA427 : full_adder port map(Sum(304), Cout(408), Sum(409), Sum(470), Cout(470));
FA428 : full_adder port map(Sum(306), Cout(409), Sum(410), Sum(471), Cout(471));
FA429 : full_adder port map(Sum(308), Cout(410), Sum(411), Sum(472), Cout(472));
FA430 : full_adder port map(Sum(310), Cout(411), Sum(412), Sum(473), Cout(473));
FA431 : full_adder port map(Sum(312), Cout(412), Sum(413), Sum(474), Cout(474));
FA432 : full_adder port map(Sum(314), Cout(413), Sum(414), Sum(475), Cout(475));
FA433 : full_adder port map(Sum(316), Cout(414), Sum(415), Sum(476), Cout(476));
FA434 : full_adder port map(Sum(318), Cout(415), Sum(416), Sum(477), Cout(477));
FA435 : full_adder port map(Sum(320), Cout(416), Sum(417), Sum(478), Cout(478));
FA436 : full_adder port map(Sum(322), Cout(417), Sum(418), Sum(479), Cout(479));
FA437 : full_adder port map(Sum(324), Cout(418), Sum(419), Sum(480), Cout(480));
FA438 : full_adder port map(Sum(326), Cout(419), Sum(420), Sum(481), Cout(481));
FA439 : full_adder port map(Sum(328), Cout(420), Sum(421), Sum(482), Cout(482));
FA440 : full_adder port map(Sum(330), Cout(421), Sum(422), Sum(483), Cout(483));
FA441 : full_adder port map(Sum(332), Cout(422), Sum(423), Sum(484), Cout(484));
FA442 : full_adder port map(Sum(334), Cout(423), Sum(424), Sum(485), Cout(485));
FA443 : full_adder port map(Sum(336), Cout(424), Sum(425), Sum(486), Cout(486));
FA444 : full_adder port map(Sum(338), Cout(425), Sum(426), Sum(487), Cout(487));
FA445 : full_adder port map(Sum(340), Cout(426), Sum(427), Sum(488), Cout(488));
FA446 : full_adder port map(Sum(342), Cout(427), Sum(428), Sum(489), Cout(489));
FA447 : full_adder port map(Sum(344), Cout(428), Sum(429), Sum(490), Cout(490));
FA448 : full_adder port map(Sum(346), Cout(429), Sum(430), Sum(491), Cout(491));
FA449 : full_adder port map(Sum(348), Cout(430), Sum(431), Sum(492), Cout(492));
FA450 : full_adder port map(Sum(350), Cout(431), Sum(432), Sum(493), Cout(493));
FA451 : full_adder port map(Sum(352), Cout(432), Sum(433), Sum(494), Cout(494));
FA452 : full_adder port map(Sum(354), Cout(433), Sum(434), Sum(495), Cout(495));
FA453 : full_adder port map(Sum(356), Cout(434), Sum(435), Sum(496), Cout(496));
FA454 : full_adder port map(Sum(358), Cout(435), Sum(436), Sum(497), Cout(497));
FA455 : full_adder port map(Sum(360), Cout(436), Sum(437), Sum(498), Cout(498));
FA456 : full_adder port map(Sum(362), Cout(437), Sum(438), Sum(499), Cout(499));
FA457 : full_adder port map(Sum(364), Cout(438), Sum(439), Sum(500), Cout(500));
FA458 : full_adder port map(Sum(366), Cout(439), Sum(440), Sum(501), Cout(501));
FA459 : full_adder port map(Sum(368), Cout(440), Sum(441), Sum(502), Cout(502));
FA460 : full_adder port map(Sum(370), Cout(441), Sum(442), Sum(503), Cout(503));
FA461 : full_adder port map(Sum(372), Cout(442), Sum(443), Sum(504), Cout(504));
FA462 : full_adder port map(Sum(374), Cout(443), Sum(444), Sum(505), Cout(505));
FA463 : full_adder port map(Sum(376), Cout(444), Sum(445), Sum(506), Cout(506));
FA464 : full_adder port map(Sum(378), Cout(445), Sum(446), Sum(507), Cout(507));
FA465 : full_adder port map(Sum(380), Cout(446), Sum(447), Sum(508), Cout(508));
FA466 : full_adder port map(Sum(382), Cout(447), Sum(448), Sum(509), Cout(509));
FA467 : full_adder port map(Sum(384), Cout(448), Sum(449), Sum(510), Cout(510));
FA468 : full_adder port map(Sum(386), Cout(449), Sum(450), Sum(511), Cout(511));
FA469 : full_adder port map(Sum(388), Cout(450), Sum(451), Sum(512), Cout(512));
FA470 : full_adder port map(Sum(390), Cout(451), Sum(452), Sum(513), Cout(513));
FA471 : full_adder port map(Sum(392), Cout(452), Sum(453), Sum(514), Cout(514));
FA472 : full_adder port map(Sum(394), Cout(453), Sum(454), Sum(515), Cout(515));
FA473 : full_adder port map(Sum(396), Cout(454), Sum(455), Sum(516), Cout(516));
FA474 : full_adder port map(Sum(398), Cout(455), Sum(456), Sum(517), Cout(517));
FA475 : full_adder port map(Sum(400), Cout(456), Sum(457), Sum(518), Cout(518));
FA476 : full_adder port map(Sum(401), Cout(457), Sum(458), Sum(519), Cout(519));
FA477 : full_adder port map(Sum(402), Cout(458), Sum(459), Sum(520), Cout(520));
FA478 : full_adder port map(Cout(402), Cout(459), Sum(460), Sum(521), Cout(521));
FA479 : full_adder port map(P(16)(30), Cout(460), Sum(461), Sum(522), Cout(522));
FA480 : full_adder port map(nSig(15), P(16)(31), Cout(461), Sum(523), Cout(523));
HA45 : half_adder port map(Sig(0), P(0)(0), Sum(524), Cout(524));
HA46 : half_adder port map(P(0)(1), Cout(524), Sum(525), Cout(525));
FA481 : full_adder port map(P(0)(2), Sum(462), Cout(525), Sum(526), Cout(526));
FA482 : full_adder port map(Cout(462), Sum(463), Cout(526), Sum(527), Cout(527));
FA483 : full_adder port map(Cout(463), Sum(464), Cout(527), Sum(528), Cout(528));
FA484 : full_adder port map(Cout(464), Sum(465), Cout(528), Sum(529), Cout(529));
FA485 : full_adder port map(Cout(465), Sum(466), Cout(529), Sum(530), Cout(530));
FA486 : full_adder port map(Cout(466), Sum(467), Cout(530), Sum(531), Cout(531));
FA487 : full_adder port map(Cout(467), Sum(468), Cout(531), Sum(532), Cout(532));
FA488 : full_adder port map(Cout(468), Sum(469), Cout(532), Sum(533), Cout(533));
FA489 : full_adder port map(Cout(469), Sum(470), Cout(533), Sum(534), Cout(534));
FA490 : full_adder port map(Cout(470), Sum(471), Cout(534), Sum(535), Cout(535));
FA491 : full_adder port map(Cout(471), Sum(472), Cout(535), Sum(536), Cout(536));
FA492 : full_adder port map(Cout(472), Sum(473), Cout(536), Sum(537), Cout(537));
FA493 : full_adder port map(Cout(473), Sum(474), Cout(537), Sum(538), Cout(538));
FA494 : full_adder port map(Cout(474), Sum(475), Cout(538), Sum(539), Cout(539));
FA495 : full_adder port map(Cout(475), Sum(476), Cout(539), Sum(540), Cout(540));
FA496 : full_adder port map(Cout(476), Sum(477), Cout(540), Sum(541), Cout(541));
FA497 : full_adder port map(Cout(477), Sum(478), Cout(541), Sum(542), Cout(542));
FA498 : full_adder port map(Cout(478), Sum(479), Cout(542), Sum(543), Cout(543));
FA499 : full_adder port map(Cout(479), Sum(480), Cout(543), Sum(544), Cout(544));
FA500 : full_adder port map(Cout(480), Sum(481), Cout(544), Sum(545), Cout(545));
FA501 : full_adder port map(Cout(481), Sum(482), Cout(545), Sum(546), Cout(546));
FA502 : full_adder port map(Cout(482), Sum(483), Cout(546), Sum(547), Cout(547));
FA503 : full_adder port map(Cout(483), Sum(484), Cout(547), Sum(548), Cout(548));
FA504 : full_adder port map(Cout(484), Sum(485), Cout(548), Sum(549), Cout(549));
FA505 : full_adder port map(Cout(485), Sum(486), Cout(549), Sum(550), Cout(550));
FA506 : full_adder port map(Cout(486), Sum(487), Cout(550), Sum(551), Cout(551));
FA507 : full_adder port map(Cout(487), Sum(488), Cout(551), Sum(552), Cout(552));
FA508 : full_adder port map(Cout(488), Sum(489), Cout(552), Sum(553), Cout(553));
FA509 : full_adder port map(Cout(489), Sum(490), Cout(553), Sum(554), Cout(554));
FA510 : full_adder port map(Cout(490), Sum(491), Cout(554), Sum(555), Cout(555));
FA511 : full_adder port map(Cout(491), Sum(492), Cout(555), Sum(556), Cout(556));
FA512 : full_adder port map(Cout(492), Sum(493), Cout(556), Sum(557), Cout(557));
FA513 : full_adder port map(Cout(493), Sum(494), Cout(557), Sum(558), Cout(558));
FA514 : full_adder port map(Cout(494), Sum(495), Cout(558), Sum(559), Cout(559));
FA515 : full_adder port map(Cout(495), Sum(496), Cout(559), Sum(560), Cout(560));
FA516 : full_adder port map(Cout(496), Sum(497), Cout(560), Sum(561), Cout(561));
FA517 : full_adder port map(Cout(497), Sum(498), Cout(561), Sum(562), Cout(562));
FA518 : full_adder port map(Cout(498), Sum(499), Cout(562), Sum(563), Cout(563));
FA519 : full_adder port map(Cout(499), Sum(500), Cout(563), Sum(564), Cout(564));
FA520 : full_adder port map(Cout(500), Sum(501), Cout(564), Sum(565), Cout(565));
FA521 : full_adder port map(Cout(501), Sum(502), Cout(565), Sum(566), Cout(566));
FA522 : full_adder port map(Cout(502), Sum(503), Cout(566), Sum(567), Cout(567));
FA523 : full_adder port map(Cout(503), Sum(504), Cout(567), Sum(568), Cout(568));
FA524 : full_adder port map(Cout(504), Sum(505), Cout(568), Sum(569), Cout(569));
FA525 : full_adder port map(Cout(505), Sum(506), Cout(569), Sum(570), Cout(570));
FA526 : full_adder port map(Cout(506), Sum(507), Cout(570), Sum(571), Cout(571));
FA527 : full_adder port map(Cout(507), Sum(508), Cout(571), Sum(572), Cout(572));
FA528 : full_adder port map(Cout(508), Sum(509), Cout(572), Sum(573), Cout(573));
FA529 : full_adder port map(Cout(509), Sum(510), Cout(573), Sum(574), Cout(574));
FA530 : full_adder port map(Cout(510), Sum(511), Cout(574), Sum(575), Cout(575));
FA531 : full_adder port map(Cout(511), Sum(512), Cout(575), Sum(576), Cout(576));
FA532 : full_adder port map(Cout(512), Sum(513), Cout(576), Sum(577), Cout(577));
FA533 : full_adder port map(Cout(513), Sum(514), Cout(577), Sum(578), Cout(578));
FA534 : full_adder port map(Cout(514), Sum(515), Cout(578), Sum(579), Cout(579));
FA535 : full_adder port map(Cout(515), Sum(516), Cout(579), Sum(580), Cout(580));
FA536 : full_adder port map(Cout(516), Sum(517), Cout(580), Sum(581), Cout(581));
FA537 : full_adder port map(Cout(517), Sum(518), Cout(581), Sum(582), Cout(582));
FA538 : full_adder port map(Cout(518), Sum(519), Cout(582), Sum(583), Cout(583));
FA539 : full_adder port map(Cout(519), Sum(520), Cout(583), Sum(584), Cout(584));
FA540 : full_adder port map(Cout(520), Sum(521), Cout(584), Sum(585), Cout(585));
FA541 : full_adder port map(Cout(521), Sum(522), Cout(585), Sum(586), Cout(586));
FA542 : full_adder port map(Cout(522), Sum(523), Cout(586), Sum(587), Cout(587));
HA47 : half_adder port map(Cout(523), Cout(587), Sum(588), Cout(588));

F1: for i in 0 to Sig'length-1 generate
	nSig(i) <= not Sig(i);
end generate;

z(0) <= Sum(524);
z(1) <= Sum(525);
z(2) <= Sum(526);
z(3) <= Sum(527);
z(4) <= Sum(528);
z(5) <= Sum(529);
z(6) <= Sum(530);
z(7) <= Sum(531);
z(8) <= Sum(532);
z(9) <= Sum(533);
z(10) <= Sum(534);
z(11) <= Sum(535);
z(12) <= Sum(536);
z(13) <= Sum(537);
z(14) <= Sum(538);
z(15) <= Sum(539);
z(16) <= Sum(540);
z(17) <= Sum(541);
z(18) <= Sum(542);
z(19) <= Sum(543);
z(20) <= Sum(544);
z(21) <= Sum(545);
z(22) <= Sum(546);
z(23) <= Sum(547);
z(24) <= Sum(548);
z(25) <= Sum(549);
z(26) <= Sum(550);
z(27) <= Sum(551);
z(28) <= Sum(552);
z(29) <= Sum(553);
z(30) <= Sum(554);
z(31) <= Sum(555);
z(32) <= Sum(556);
z(33) <= Sum(557);
z(34) <= Sum(558);
z(35) <= Sum(559);
z(36) <= Sum(560);
z(37) <= Sum(561);
z(38) <= Sum(562);
z(39) <= Sum(563);
z(40) <= Sum(564);
z(41) <= Sum(565);
z(42) <= Sum(566);
z(43) <= Sum(567);
z(44) <= Sum(568);
z(45) <= Sum(569);
z(46) <= Sum(570);
z(47) <= Sum(571);
z(48) <= Sum(572);
z(49) <= Sum(573);
z(50) <= Sum(574);
z(51) <= Sum(575);
z(52) <= Sum(576);
z(53) <= Sum(577);
z(54) <= Sum(578);
z(55) <= Sum(579);
z(56) <= Sum(580);
z(57) <= Sum(581);
z(58) <= Sum(582);
z(59) <= Sum(583);
z(60) <= Sum(584);
z(61) <= Sum(585);
z(62) <= Sum(586);
z(63) <= Sum(587);

end architecture;