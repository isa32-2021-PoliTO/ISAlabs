package const_MEM is

   constant ADDRESS_LENGTH : natural := 16;
   constant DATA_LENGTH : natural := 32;

end const_MEM;
